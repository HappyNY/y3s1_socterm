module GPPCU_INSTR_DEC #(
    
)
(
    
);
    
    

endmodule