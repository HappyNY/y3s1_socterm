module GPPCU_STALL_GEN(
    
);


endmodule